`define AE0_PRESENT 1
//`define AE1_PRESENT 1
//`define AE2_PRESENT 1
//`define AE3_PRESENT 1
